library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
library work;

ENTITY testbench_phase2 IS
END testbench_phase2;

ARCHITECTURE testbench_arch OF testbench_phase2 IS

signal ren0_tb   		;  
signal ren1_tb   		;  
signal ren2_tb   		;  
signal ren3_tb   		;  
signal ren4_tb   		;  
signal ren5_tb   		;  
signal ren6_tb   		;  
signal ren7_tb   		;  
signal ren8_tb   		;  
signal ren9_tb   		;  
signal renA_tb   		;  
signal renB_tb   		;  
signal renC_tb   		;  
signal renD_tb   		;  
signal renE_tb   		;  
signal renF_tb   		;  
signal   clr_tb  		;    
signal   clk_tb  		;    
signal R0out_tb  		;  
signal R1out_tb  		;  
signal R2out_tb  		;  
signal R3out_tb  		;  
signal R4out_tb  		;  
signal R5out_tb  		;  
signal R6out_tb  		;  
signal R7out_tb  		;  
signal R8out_tb  		;  
signal R9out_tb  		;  
signal R10out_tb 		;  
signal R11out_tb 		;  
signal R12out_tb 		;  
signal R13out_tb 		;  
signal R14out_tb 		;  
signal R15out_tb 		;  
signal Zhighout_tb 	;
signal Zlowout_tb  	;
signal InPortout_tb	;
signal HIin_tb     	;
signal PCin_tb     	;
signal LOin_tb     	;
signal MDRin_tb    	;
signal HIoutEn_tb  	;
signal LOoutEn_tb  	;
signal PCoutEn_tb  	;
signal MDRoutEn_tb 	;
signal CoutEn_tb 		; 
signal reny_tb			; 	  
signal renz_tb			; 	  
signal ReadIn_tb		; 	  
signal WriteEn_tb		;    
signal MARin_tb		;  	  
signal IRen_tb			;  	  
signal CONin_tb		;  	  
signal OUTen_tb		;  	  
signal Strobe_tb		;  	  
signal Gra_tb			;  	  
signal Grb_tb			;  	  
signal Grc_tb			;  	  
signal SelEncin_tb	;   
signal SelEncout_tb	;  
signal BAout_tb		;  	  
signal Empty_tb		; 	  
signal HIout_tb		;  	  
signal InPortIn_tb	;   
signal LOout_tb		;  	  
signal Mdatain_tb		;    
signal MDRout_tb		;  	  
signal operation_tb	;  
signal PCout_tb		;      
signal rout0_tb		;      
signal rout1_tb		;      
signal rout2_tb		;      
signal rout3_tb		;      
signal rout4_tb		;      
signal rout5_tb		;      
signal rout6_tb		;      
signal rout7_tb		;      
signal rout8_tb		;      
signal rout9_tb		;      
signal routa_tb		;      
signal routb_tb		;      
signal routc_tb		;      
signal routd_tb		;      
signal route_tb		;      
signal routf_tb		;      
signal routy_tb		;      
signal Zhigh_tb		;      
signal Zlow_tb			;       
signal CONout_tb		;  	  
signal Address_tb		; 	  
signal IRout_tb		;  	  
signal Out_Port_tb	;   
signal RALLin_tb		;  	  
signal RALLout_tb		;    


component ELEC374 
PORT
	(
		ren0 :  IN  STD_LOGIC;
		ren1 :  IN  STD_LOGIC;
		ren2 :  IN  STD_LOGIC;
		ren3 :  IN  STD_LOGIC;
		ren4 :  IN  STD_LOGIC;
		ren5 :  IN  STD_LOGIC;
		ren6 :  IN  STD_LOGIC;
		ren7 :  IN  STD_LOGIC;
		ren8 :  IN  STD_LOGIC;
		ren9 :  IN  STD_LOGIC;
		renA :  IN  STD_LOGIC;
		renB :  IN  STD_LOGIC;
		renC :  IN  STD_LOGIC;
		renD :  IN  STD_LOGIC;
		renE :  IN  STD_LOGIC;
		renF :  IN  STD_LOGIC;
		clr :  IN  STD_LOGIC;
		clk :  IN  STD_LOGIC;
		R0out :  IN  STD_LOGIC;
		R1out :  IN  STD_LOGIC;
		R2out :  IN  STD_LOGIC;
		R3out :  IN  STD_LOGIC;
		R4out :  IN  STD_LOGIC;
		R5out :  IN  STD_LOGIC;
		R6out :  IN  STD_LOGIC;
		R7out :  IN  STD_LOGIC;
		R8out :  IN  STD_LOGIC;
		R9out :  IN  STD_LOGIC;
		R10out :  IN  STD_LOGIC;
		R11out :  IN  STD_LOGIC;
		R12out :  IN  STD_LOGIC;
		R13out :  IN  STD_LOGIC;
		R14out :  IN  STD_LOGIC;
		R15out :  IN  STD_LOGIC;
		Zhighout :  IN  STD_LOGIC;
		Zlowout :  IN  STD_LOGIC;
		InPortout :  IN  STD_LOGIC;
		HIin :  IN  STD_LOGIC;
		PCin :  IN  STD_LOGIC;
		LOin :  IN  STD_LOGIC;
		MDRin :  IN  STD_LOGIC;
		HIoutEn :  IN  STD_LOGIC;
		LOoutEn :  IN  STD_LOGIC;
		PCoutEn :  IN  STD_LOGIC;
		MDRoutEn :  IN  STD_LOGIC;
		CoutEn :  IN  STD_LOGIC;
		reny :  IN  STD_LOGIC;
		renz :  IN  STD_LOGIC;
		ReadIn :  IN  STD_LOGIC;
		WriteEn :  IN  	STD_LOGIC;
		MARin :  IN  		STD_LOGIC;
		IRen :  IN  		STD_LOGIC;
		CONin :  IN  		STD_LOGIC;
		OUTen :  IN  		STD_LOGIC;
		Strobe :  IN  		STD_LOGIC;
		Gra :  IN  			STD_LOGIC;
		Grb :  IN  			STD_LOGIC;
		Grc :  IN  			STD_LOGIC;
		SelEncin :  IN  	STD_LOGIC;
		SelEncout :  IN  	STD_LOGIC;
		BAout :  IN  		STD_LOGIC;
		Empty :  IN  		STD_LOGIC_VECTOR(31 DOWNTO 0);
		HIout :  INOUT  	STD_LOGIC_VECTOR(31 DOWNTO 0);
		InPortIn :  IN  	STD_LOGIC_VECTOR(31 DOWNTO 0);
		LOout :  INOUT  	STD_LOGIC_VECTOR(31 DOWNTO 0);
		Mdatain :  IN  	STD_LOGIC_VECTOR(31 DOWNTO 0);
		MDRout :  INOUT  	STD_LOGIC_VECTOR(31 DOWNTO 0);
		operation :  IN  	STD_LOGIC_VECTOR(3 DOWNTO 0);
		PCout :  INOUT  	STD_LOGIC_VECTOR(31 DOWNTO 0);
		rout0 :  INOUT  	STD_LOGIC_VECTOR(31 DOWNTO 0);
		rout1 :  INOUT  	STD_LOGIC_VECTOR(31 DOWNTO 0);
		rout2 :  INOUT  	STD_LOGIC_VECTOR(31 DOWNTO 0);
		rout3 :  INOUT  	STD_LOGIC_VECTOR(31 DOWNTO 0);
		rout4 :  INOUT  	STD_LOGIC_VECTOR(31 DOWNTO 0);
		rout5 :  INOUT  	STD_LOGIC_VECTOR(31 DOWNTO 0);
		rout6 :  INOUT  	STD_LOGIC_VECTOR(31 DOWNTO 0);
		rout7 :  INOUT  	STD_LOGIC_VECTOR(31 DOWNTO 0);
		rout8 :  INOUT  	STD_LOGIC_VECTOR(31 DOWNTO 0);
		rout9 :  INOUT  	STD_LOGIC_VECTOR(31 DOWNTO 0);
		routa :  INOUT  	STD_LOGIC_VECTOR(31 DOWNTO 0);
		routb :  INOUT  	STD_LOGIC_VECTOR(31 DOWNTO 0);
		routc :  INOUT  	STD_LOGIC_VECTOR(31 DOWNTO 0);
		routd :  INOUT  	STD_LOGIC_VECTOR(31 DOWNTO 0);
		route :  INOUT  	STD_LOGIC_VECTOR(31 DOWNTO 0);
		routf :  INOUT  	STD_LOGIC_VECTOR(31 DOWNTO 0);
		routy :  INOUT  	STD_LOGIC_VECTOR(31 DOWNTO 0);
		Zhigh :  INOUT  	STD_LOGIC_VECTOR(31 DOWNTO 0);
		Zlow :  INOUT 		STD_LOGIC_VECTOR(31 DOWNTO 0);
		CONout :  OUT 		STD_LOGIC;
		Address :  OUT  	STD_LOGIC_VECTOR(8 DOWNTO 0);
		IRout :  OUT  		STD_LOGIC_VECTOR(31 DOWNTO 0);
		Out_Port :  OUT  	STD_LOGIC_VECTOR(31 DOWNTO 0);
		RALLin :  OUT  	STD_LOGIC_VECTOR(15 DOWNTO 0);
		RALLout :  OUT  	STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
	end component ELEC374;
	
	
end architecture testbench_arch;